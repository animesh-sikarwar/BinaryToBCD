`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module bin_2_7seg(input [3:0] a , output reg [6:0] b

    );
    always @(a)
    case(a) 
    4'd0:b=7'b1111110;
    4'd1:b=7'b0110000;
    4'd2:b=7'b1101101;
    4'd3:b=7'b1111001;
    4'd4:b=7'b0110011;
    4'd5:b=7'b1011011;
    4'd6:b=7'b1011111;
    4'd7:b=7'b1110000;
    4'd8:b=7'b1111111;
    4'd9:b=7'b1111011;
    default:b=7'b0000000;
    endcase
    
    
endmodule
